//==============================================================
// File        : fetch.v
// Description : Instruction memory + PC logic
// Author      : Mauro Ferreira
//==============================================================

module fetch (
    input clk, rst,
    output reg [31:0] pc,
    output [31:0] instruction
);

    // Simple instruction memory with 256 32-bit instructions
    reg [31:0] instr_mem [0:255];

    // Instruction 32 bit set
	initial begin
    instr_mem[0]  = 32'b0000000_00010_00001_000_00011_0110011; // ADD x3, x1, x2
    instr_mem[1]  = 32'b0100000_00011_00010_000_00100_0110011; // SUB x4, x2, x3
    instr_mem[2]  = 32'b0000000_00100_00011_111_00101_0110011; // AND x5, x3, x4
    instr_mem[3]  = 32'b0000000_00101_00100_110_00110_0110011; // OR  x6, x4, x5
    instr_mem[4]  = 32'b0000000_00110_00101_100_00111_0110011; // XOR x7, x5, x6
    instr_mem[5]  = 32'b0000000_00001_00001_000_00001_0110011; // ADD x1, x1, x1
    instr_mem[6]  = 32'b0000000_00010_00010_000_00010_0110011; // ADD x2, x2, x2
    instr_mem[7]  = 32'b0000000_00011_00011_000_00011_0110011; // ADD x3, x3, x3
    instr_mem[8]  = 32'b0100000_00011_00001_000_00100_0110011; // SUB x4, x1, x3
    instr_mem[9]  = 32'b0000000_00010_00011_000_00101_0110011; // ADD x5, x3, x2
    instr_mem[10] = 32'b0100000_00010_00001_000_00110_0110011; // SUB x6, x1, x2
    instr_mem[11] = 32'b0000000_00001_00010_111_00111_0110011; // AND x7, x2, x1
    instr_mem[12] = 32'b0000000_00111_00110_110_00001_0110011; // OR  x1, x6, x7
    instr_mem[13] = 32'b0000000_00101_00100_100_00010_0110011; // XOR x2, x4, x5
    instr_mem[14] = 32'b0000000_00100_00001_000_00011_0110011; // ADD x3, x1, x4
    instr_mem[15] = 32'b0000000_00111_00101_000_00100_0110011; // ADD x4, x5, x7
    instr_mem[16] = 32'b0100000_00010_00011_000_00101_0110011; // SUB x5, x3, x2
    instr_mem[17] = 32'b0000000_00001_00011_111_00110_0110011; // AND x6, x3, x1
    instr_mem[18] = 32'b0000000_00010_00100_110_00111_0110011; // OR  x7, x4, x2
    instr_mem[19] = 32'b0000000_00110_00010_100_00001_0110011; // XOR x1, x2, x6
    instr_mem[20] = 32'b0000000_00100_00110_000_00010_0110011; // ADD x2, x6, x4
    instr_mem[21] = 32'b0100000_00101_00100_000_00011_0110011; // SUB x3, x4, x5
    instr_mem[22] = 32'b0000000_00101_00011_111_00100_0110011; // AND x4, x3, x5
    instr_mem[23] = 32'b0000000_00010_00011_110_00101_0110011; // OR  x5, x3, x2
    instr_mem[24] = 32'b0000000_00100_00111_100_00110_0110011; // XOR x6, x7, x4
    instr_mem[25] = 32'b0000000_00001_00001_000_00001_0110011; // ADD x1, x1, x1
    instr_mem[26] = 32'b0000000_00010_00010_000_00010_0110011; // ADD x2, x2, x2
    instr_mem[27] = 32'b0000000_00011_00011_000_00011_0110011; // ADD x3, x3, x3
    instr_mem[28] = 32'b0100000_00011_00001_000_00100_0110011; // SUB x4, x1, x3
    instr_mem[29] = 32'b0000000_00010_00011_000_00101_0110011; // ADD x5, x3, x2
    instr_mem[30] = 32'b0000000_00001_00010_111_00110_0110011; // AND x6, x2, x1
    instr_mem[31] = 32'b0000000_00111_00110_110_00111_0110011; // OR  x7, x6, x7
	end
    assign instruction = instr_mem[pc >> 2]; // Word-aligned access

    always @(posedge clk or posedge rst) begin
        if (rst)
            pc <= 0;
        else
            pc <= pc + 4; // Advance to next instruction
    end

endmodule
